-- Top level entity, MARK_II SoC
--
-- Part of MARK II project. For informations about license, please
-- see file /LICENSE .
--
-- author: Vladislav Mlejnecký
-- email: v.mlejnecky@seznam.cz

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MARK_II is
    port(
        --control signals
        clk: in std_logic;
        res: in std_logic;

        --gpio
        porta: inout std_logic_vector(7 downto 0);
        portb: inout std_logic_vector(7 downto 0);

        --timers
        tim0_pwma: out std_logic;
        tim0_pwmb: out std_logic;
        tim1_pwma: out std_logic;
        tim1_pwmb: out std_logic;
        tim2_pwma: out std_logic;
        tim2_pwmb: out std_logic;
        tim3_pwma: out std_logic;
        tim3_pwmb: out std_logic;

        --uarts
        tx0: out std_logic;
        rx0: in std_logic;
        tx1: out std_logic;
        rx1: in std_logic;
        tx2: out std_logic;
        rx2: in std_logic;

        --vga
        h_sync: out std_logic;
        v_sync: out std_logic;
        red: out std_logic_vector(1 downto 0);
        green: out std_logic_vector(1 downto 0);
        blue: out std_logic_vector(1 downto 0);

        --keyboard
        ps2clk: in std_logic;
        ps2dat: in std_logic
    );
end entity MARK_II;

architecture MARK_II_arch of MARK_II is

    attribute chip_pin : string;

    attribute chip_pin of clk           : signal is "R8";
    attribute chip_pin of res           : signal is "J15";

    attribute chip_pin of porta         : signal is "L3, B1, F3, D1, A11, B13, A13, A15";
    attribute chip_pin of portb         : signal is "A2, A3, B3, B4, A4, B5, A5, D5";

    attribute chip_pin of tim0_pwma     : signal is "B6";
    attribute chip_pin of tim0_pwmb     : signal is "A6";
    attribute chip_pin of tim1_pwma     : signal is "B7";
    attribute chip_pin of tim1_pwmb     : signal is "D6";
    attribute chip_pin of tim2_pwma     : signal is "A7";
    attribute chip_pin of tim2_pwmb     : signal is "C6";
    attribute chip_pin of tim3_pwma     : signal is "C8";
    attribute chip_pin of tim3_pwmb     : signal is "E6";

    attribute chip_pin of tx0           : signal is "J16";
    attribute chip_pin of rx0           : signal is "J13";
    attribute chip_pin of tx1           : signal is "K15";
    attribute chip_pin of rx1           : signal is "N14";
    attribute chip_pin of tx2           : signal is "E11";
    attribute chip_pin of rx2           : signal is "E10";

    attribute chip_pin of h_sync        : signal is "L14";
    attribute chip_pin of v_sync        : signal is "M10";
    attribute chip_pin of red           : signal is "N15,R14";
    attribute chip_pin of green         : signal is "N16,P15";
    attribute chip_pin of blue          : signal is "P16,R16";

    attribute chip_pin of ps2clk        : signal is "L16";
    attribute chip_pin of ps2dat        : signal is "L15";

    component cpu is
        port(
            --system interface
            clk: in std_logic;
            res: in std_logic;
            --bus interface
            address: out std_logic_vector(23 downto 0);
            data_mosi: out std_logic_vector(31 downto 0);
            data_miso: in std_logic_vector(31 downto 0);
            we: out std_logic;
            oe: out std_logic;
            ack: in std_logic;
            swirq: out std_logic;
            --interrupts
            int: in std_logic;
            int_address: in std_logic_vector(23 downto 0);
            int_accept: out std_logic;
            int_completed: out std_logic
        );
    end component cpu;

    component intController is
        generic(
            BASE_ADDRESS: unsigned(23 downto 0) := x"000000"    --base address
        );
        port(
            --bus
            clk: in std_logic;
            res: in std_logic;
            address: in std_logic_vector(23 downto 0);
            data_mosi: in std_logic_vector(31 downto 0);
            data_miso: out std_logic_vector(31 downto 0);
            WR: in std_logic;
            RD: in std_logic;
            ack: out std_logic;
            --device
            int_req: in std_logic_vector(15 downto 0);      --peripherals may request interrupt with this signal
            int_accept: in std_logic;                       --from the CPU
            int_completed: in std_logic;                    --from the CPU
            int_cpu_address: out std_logic_vector(23 downto 0);  --connect this to the CPU, this is address of ISR
            int_cpu_rq: out std_logic
        );
    end component intController;

    component gpio is
        generic(
            BASE_ADDRESS: unsigned(23 downto 0) := x"000000";    --base address of the GPIO
            GPIO_WIDE: natural := 32       --wide of the gpios
        );
        port(
            clk: in std_logic;
            res: in std_logic;
            address: in std_logic_vector(23 downto 0);
            data_mosi: in std_logic_vector(31 downto 0);
            data_miso: out std_logic_vector(31 downto 0);
            WR: in std_logic;
            RD: in std_logic;
            ack: out std_logic;
            --outputs
            port_a: inout std_logic_vector((GPIO_WIDE-1) downto 0);
            port_b: inout std_logic_vector((GPIO_WIDE-1) downto 0)
        );
    end component gpio;

    component rom is
        generic(
            BASE_ADDRESS: unsigned(23 downto 0) := x"000000"    --base address of the ROM
        );
        port(
            clk: in std_logic;
            res: in std_logic;
            address: in std_logic_vector(23 downto 0);
            data_mosi: in std_logic_vector(31 downto 0);
            data_miso: out std_logic_vector(31 downto 0);
            WR: in std_logic;
            RD: in std_logic;
            ack: out std_logic
        );
    end component rom;

    component ram is
        generic(
            BASE_ADDRESS: unsigned(23 downto 0) := x"000000";    --base address of the RAM
            ADDRESS_WIDE: natural := 8  --default address range
        );
        port(
            clk: in std_logic;
            res: in std_logic;
            address: in std_logic_vector(23 downto 0);
            data_mosi: in std_logic_vector(31 downto 0);
            data_miso: out std_logic_vector(31 downto 0);
            WR: in std_logic;
            RD: in std_logic;
            ack: out std_logic
        );
    end component ram;

    component systim is
        generic(
            BASE_ADDRESS: unsigned(23 downto 0) := x"000000"    --base address
        );
        port(
            --bus
            clk: in std_logic;
            res: in std_logic;
            address: in std_logic_vector(23 downto 0);
            data_mosi: in std_logic_vector(31 downto 0);
            data_miso: out std_logic_vector(31 downto 0);
            WR: in std_logic;
            RD: in std_logic;
            ack: out std_logic;
            --device
            intrq: out std_logic
        );
    end component systim;

    component timer is
        generic(
            BASE_ADDRESS: unsigned(23 downto 0) := x"000000"    --base address
        );
        port(
            --bus
            clk: in std_logic;
            res: in std_logic;
            address: in std_logic_vector(23 downto 0);
            data_mosi: in std_logic_vector(31 downto 0);
            data_miso: out std_logic_vector(31 downto 0);
            WR: in std_logic;
            RD: in std_logic;
            ack: out std_logic;
            --device
            pwma: out std_logic;
            pwmb: out std_logic;
            intrq: out std_logic
        );
    end component;

    component uart is
        generic(
            BASE_ADDRESS: unsigned(23 downto 0) := x"000000"    --base address of the GPIO
        );
        port(
            clk: in std_logic;
            res: in std_logic;
            address: in std_logic_vector(23 downto 0);
            data_mosi: in std_logic_vector(31 downto 0);
            data_miso: out std_logic_vector(31 downto 0);
            WR: in std_logic;
            RD: in std_logic;
            ack: out std_logic;
            --device
            clk_uart: in std_logic;
            rx: in std_logic;
            tx: out std_logic;
            intrq: out std_logic
        );
    end component uart;

    component vga is
        generic(
            BASE_ADDRESS: unsigned(23 downto 0) := x"000000"    --base address of the RAM
        );
        port(
            clk_bus: in std_logic;
            address: in std_logic_vector(23 downto 0);
            data_mosi: in std_logic_vector(31 downto 0);
            data_miso: out std_logic_vector(31 downto 0);
            WR: in std_logic;
            RD: in std_logic;
            ack: out std_logic;
            --device
            clk_31M5: in std_logic;
            h_sync: out std_logic;
            v_sync: out std_logic;
            red: out std_logic_vector(1 downto 0);
            green: out std_logic_vector(1 downto 0);
            blue: out std_logic_vector(1 downto 0)
        );
    end component vga;

    component ps2 is
        generic(
            BASE_ADDRESS: unsigned(23 downto 0) := x"000000"
        );
        port(
            clk: in std_logic;
            res: in std_logic;
            address: in std_logic_vector(23 downto 0);
            data_miso: out std_logic_vector(31 downto 0);
            RD: in std_logic;
            ack: out std_logic;
            --device
            ps2clk: in std_logic;
            ps2dat: in std_logic;
            intrq: out std_logic
        );
    end component ps2;

    component pll
        port(
            inclk0: in std_logic:= '0';
            c0: out std_logic;
            c1: out std_logic;
            c2: out std_logic
        );
    end component;

    --signal for internal bus
    signal bus_address: std_logic_vector(23 downto 0);
    signal bus_data_mosi, bus_data_miso: std_logic_vector(31 downto 0);
    signal bus_ack, bus_WR, bus_RD: std_logic;
    signal int_req: std_logic_vector(15 downto 0) := x"0000";

    --signal for interconnect CPU and int controller
    signal intCompleted, intAccepted: std_logic;
    signal intCPUReq: std_logic;
    signal intAddress: std_logic_vector(23 downto 0);

    signal clk_31M5: std_logic;     -- 31,5 MHz clk for vga
    signal clk_uart: std_logic;     -- 14,4 MHz clk for uarts
    signal clk_sys: std_logic;      -- 50 MHz clk for CPU

    signal resi: std_logic;         --inverted reset

    signal rom_ack, ram_ack, int_ack, gpio_ack, systim_ack, vga_ack, tim0_ack, ram1_ack,
           tim1_ack,tim2_ack,tim3_ack, uart0_ack, uart1_ack, uart2_ack, ps2_ack : std_logic;

begin

    resi <= not(res);
   
    pll0: pll
        port map(clk, clk_uart, clk_31M5, clk_sys);
    
    cpu0: cpu
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, bus_ack, int_req(0), intCPUReq, intAddress, intAccepted, intCompleted);

    int0: intController
        generic map(x"00010F")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, int_ack, int_req, intAccepted, intCompleted, intAddress, intCPUReq);

    systim0: systim
        generic map(x"000104")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, systim_ack, int_req(1));

    gpio0: gpio
        generic map(x"000100", 8)
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, gpio_ack, porta, portb);

    rom0: rom
        generic map(x"000000")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, rom_ack);

    ram0: ram
        generic map(x"000400", 10)
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, ram_ack);

    tim0: timer
        generic map(x"000120")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, tim0_ack, tim0_pwma, tim0_pwmb, int_req(12));

    tim1: timer
        generic map(x"000124")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, tim1_ack, tim1_pwma, tim1_pwmb, int_req(13));

    tim2: timer
        generic map(x"000128")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, tim2_ack, tim2_pwma, tim2_pwmb, int_req(14));

    tim3: timer
        generic map(x"00012C")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, tim3_ack, tim3_pwma, tim3_pwmb, int_req(15));

    uart0: uart
        generic map(x"000130")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, uart0_ack, clk_uart, rx0, tx0, int_req(8));

    uart1: uart
        generic map(x"000134")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, uart1_ack, clk_uart, rx1, tx1, int_req(9));

    uart2: uart
        generic map(x"000138")
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, uart2_ack, clk_uart, rx2, tx2, int_req(10));

    vga0: vga
        generic map(x"001000")
        port map(clk_sys, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, vga_ack, clk_31M5, h_sync, v_sync, red, green, blue);

    ps2keyboard0: ps2
        generic map(x"000106")
        port map(clk_sys, resi, bus_address, bus_data_miso, bus_RD, ps2_ack, ps2clk, ps2dat, int_req(11));

    ram1: ram
        generic map(x"100000", 13)
        port map(clk_sys, resi, bus_address, bus_data_mosi, bus_data_miso, bus_WR, bus_RD, ram1_ack);

    bus_ack <=
        rom_ack or ram_ack or int_ack or gpio_ack or systim_ack or vga_ack or tim0_ack or
        tim1_ack or tim2_ack or tim3_ack or uart0_ack or uart1_ack or uart2_ack or ps2_ack or ram1_ack;

end architecture MARK_II_arch;
