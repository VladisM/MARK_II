-- Read only memory with font.
--
-- Part of MARK_II SoC project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity font_rom is
    port(
        clk: in std_logic;
        addr: in unsigned(10 downto 0);
        data: out unsigned(7 downto 0)
    );
end entity font_rom;

architecture font_rom_arch of font_rom is

    type rom_type is array (0 to 2**11-1) of unsigned(7 downto 0);

    constant ROM: rom_type :=(
        -- code 0x00
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        -- code 0x01
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "11111111",
        "11111111",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x02
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "11111111",
        "11111111",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        -- code 0x03
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "11111000",
        "11111000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        -- code 0x04
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011111",
        "00011111",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        -- code 0x05
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "11111000",
        "11111000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x06
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011111",
        "00011111",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x07
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011111",
        "00011111",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        -- code 0x08
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "11111000",
        "11111000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        -- code 0x09
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "11111111",
        "11111111",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        -- code 0x0A
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "11111111",
        "11111111",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x0B
        "00000000",
        "00000000",
        "01000000",
        "01100000",
        "01110000",
        "01111000",
        "01111100",
        "01111110",
        "01111110",
        "01111100",
        "01111000",
        "01110000",
        "01100000",
        "01000000",
        "00000000",
        "00000000",
        -- code 0x0C
        "00000000",
        "00000000",
        "00000010",
        "00000110",
        "00001110",
        "00011110",
        "00111110",
        "01111110",
        "01111110",
        "00111110",
        "00011110",
        "00001110",
        "00000110",
        "00000010",
        "00000000",
        "00000000",
        -- code 0x0D
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00011000",
        "00111100",
        "00111100",
        "00111100",
        "01111110",
        "01111110",
        "01111110",
        "11111111",
        "11111111",
        "11111111",
        "00000000",
        "00000000",
        -- code 0x0E
        "00000000",
        "00000000",
        "11111111",
        "11111111",
        "11111111",
        "01111110",
        "01111110",
        "01111110",
        "00111100",
        "00111100",
        "00111100",
        "00011000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        -- code 0x0F
        "11011011",
        "00100100",
        "11011011",
        "00100100",
        "11011011",
        "00100100",
        "11011011",
        "00100100",
        "11011011",
        "00100100",
        "11011011",
        "00100100",
        "11011011",
        "00100100",
        "11011011",
        "00100100",
        -- code 0x10
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        "11111111",
        -- code 0x11
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00110000",
        "00011000",
        "00001100",
        "01111110",
        "01111110",
        "00001100",
        "00011000",
        "00110000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x12
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00001100",
        "00011000",
        "00110000",
        "01111110",
        "01111110",
        "00110000",
        "00011000",
        "00001100",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x13
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00011000",
        "10011001",
        "11011011",
        "01111110",
        "00111100",
        "00011000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x14
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00111100",
        "01111110",
        "11011011",
        "10011001",
        "00011000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x15
        "00000000",
        "00110000",
        "01001000",
        "01001000",
        "00110000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x16
        "00000000",
        "00000000",
        "00000000",
        "01001000",
        "01001000",
        "00100100",
        "00100100",
        "00010010",
        "00010010",
        "00100100",
        "00100100",
        "01001000",
        "01001000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x17
        "00000000",
        "00000000",
        "00000000",
        "00010010",
        "00010010",
        "00100100",
        "00100100",
        "01001000",
        "01001000",
        "00100100",
        "00100100",
        "00010010",
        "00010010",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x18
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00110110",
        "01111111",
        "01111111",
        "01111111",
        "01111111",
        "00111110",
        "00011100",
        "00001000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x19
        "00000000",
        "00000000",
        "00001000",
        "00011100",
        "00011100",
        "00111110",
        "00111110",
        "01111111",
        "00111110",
        "00111110",
        "00011100",
        "00011100",
        "00001000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x1A
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00111100",
        "00111100",
        "11100111",
        "11100111",
        "11100111",
        "11100111",
        "00011000",
        "00011000",
        "00111100",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x1B
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00111100",
        "01111110",
        "11111111",
        "11111111",
        "01111110",
        "00011000",
        "00011000",
        "00111100",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x1C
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01000010",
        "01000010",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x1D
        "00000000",
        "00000000",
        "01111110",
        "01100110",
        "01111110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01101110",
        "01101110",
        "11101100",
        "11100000",
        "11000000",
        "00000000",
        "00000000",
        -- code 0x1E
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "00000000",
        "00000000",
        "00000000",
        "01000010",
        "00111100",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x1F
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "01000010",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x20
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x21
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00000000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        -- code 0x22
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x23
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "11111111",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "11111111",
        "01100110",
        "01100110",
        "01100110",
        "00000000",
        "00000000",
        -- code 0x24
        "00011000",
        "00011000",
        "00111100",
        "01100110",
        "01100010",
        "01100000",
        "01100000",
        "00111100",
        "00000110",
        "00000110",
        "00000110",
        "01000110",
        "01100110",
        "00111100",
        "00011000",
        "00011000",
        -- code 0x25
        "00000000",
        "00000000",
        "00100010",
        "01010010",
        "01010100",
        "00100100",
        "00001000",
        "00001000",
        "00010000",
        "00010000",
        "00100100",
        "00101010",
        "01001010",
        "01000100",
        "00000000",
        "00000000",
        -- code 0x26
        "00000000",
        "00000000",
        "00000000",
        "00111000",
        "01101100",
        "01101100",
        "00111000",
        "01110000",
        "11011010",
        "11001100",
        "11001100",
        "11001100",
        "11001100",
        "01110110",
        "00000000",
        "00000000",
        -- code 0x27
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x28
        "00000000",
        "00001100",
        "00011100",
        "00011000",
        "00111000",
        "00110000",
        "00110000",
        "01110000",
        "01110000",
        "00110000",
        "00110000",
        "00111000",
        "00011000",
        "00011100",
        "00001100",
        "00000000",
        -- code 0x29
        "00000000",
        "00110000",
        "00111000",
        "00011000",
        "00011100",
        "00001100",
        "00001100",
        "00001110",
        "00001110",
        "00001100",
        "00001100",
        "00011100",
        "00011000",
        "00111000",
        "00110000",
        "00000000",
        -- code 0x2A
        "00000000",
        "00000000",
        "00011000",
        "01011010",
        "00111100",
        "00111100",
        "01011010",
        "00011000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x2B
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "01111110",
        "01111110",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x2C
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00011000",
        "00110000",
        -- code 0x2D
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01111110",
        "01111110",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x2E
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        -- code 0x2F
        "00000000",
        "00000000",
        "00000010",
        "00000110",
        "00000110",
        "00001100",
        "00001100",
        "00011000",
        "00011000",
        "00110000",
        "00110000",
        "01100000",
        "01100000",
        "01000000",
        "00000000",
        "00000000",
        -- code 0x30
        "00000000",
        "00000000",
        "00011000",
        "00111100",
        "01100110",
        "01100110",
        "01110110",
        "01110110",
        "01101110",
        "01101110",
        "01100110",
        "01100110",
        "00111100",
        "00011000",
        "00000000",
        "00000000",
        -- code 0x31
        "00000000",
        "00000000",
        "00001000",
        "00011000",
        "00111000",
        "01111000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "01111110",
        "00000000",
        "00000000",
        -- code 0x32
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "00000110",
        "00000110",
        "00000110",
        "00001100",
        "00011000",
        "00110000",
        "01100000",
        "01100010",
        "01111110",
        "00000000",
        "00000000",
        -- code 0x33
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "00000110",
        "00000110",
        "00000110",
        "00111100",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x34
        "00000000",
        "00000000",
        "00001100",
        "00011100",
        "00011100",
        "00101100",
        "00101100",
        "01001100",
        "01001100",
        "01111110",
        "00001100",
        "00001100",
        "00001100",
        "00011110",
        "00000000",
        "00000000",
        -- code 0x35
        "00000000",
        "00000000",
        "01111110",
        "01100000",
        "01100000",
        "01100000",
        "01100000",
        "01111100",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x36
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100000",
        "01100000",
        "01100000",
        "01111100",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x37
        "00000000",
        "00000000",
        "01111110",
        "01100110",
        "00000110",
        "00000110",
        "00001110",
        "00001100",
        "00011100",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        -- code 0x38
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x39
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111110",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "01000110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x3A
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x3B
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00011000",
        "00110000",
        -- code 0x3C
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000100",
        "00001100",
        "00011000",
        "00110000",
        "00110000",
        "00011000",
        "00001100",
        "00000100",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x3D
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01111110",
        "01111110",
        "00000000",
        "00000000",
        "01111110",
        "01111110",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x3E
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00100000",
        "00110000",
        "00011000",
        "00001100",
        "00001100",
        "00011000",
        "00110000",
        "00100000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x3F
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "00000110",
        "00001100",
        "00011000",
        "00011000",
        "00011000",
        "00000000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        -- code 0x40
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "01101110",
        "01101110",
        "01101110",
        "01101110",
        "01101100",
        "01100000",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x41
        "00000000",
        "00000000",
        "00011000",
        "00111100",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01111110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00000000",
        "00000000",
        -- code 0x42
        "00000000",
        "00000000",
        "01111100",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "00111100",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "01111100",
        "00000000",
        "00000000",
        -- code 0x43
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100010",
        "01100000",
        "01100000",
        "01100000",
        "01100000",
        "01100000",
        "01100000",
        "01100010",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x44
        "00000000",
        "00000000",
        "01111100",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "00110010",
        "01111100",
        "00000000",
        -- code 0x45
        "00000000",
        "00000000",
        "01111110",
        "00110010",
        "00110000",
        "00110000",
        "00110000",
        "00111100",
        "00111100",
        "00110000",
        "00110000",
        "00110000",
        "00110010",
        "01111110",
        "00000000",
        "00000000",
        -- code 0x46
        "00000000",
        "00000000",
        "01111110",
        "00110010",
        "00110000",
        "00110000",
        "00110000",
        "00111100",
        "00111100",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "01111000",
        "00000000",
        "00000000",
        -- code 0x47
        "00000000",
        "00000000",
        "00111100",
        "01100010",
        "01100000",
        "01100000",
        "01100000",
        "01100000",
        "01101110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111010",
        "00000000",
        "00000000",
        -- code 0x48
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01111110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00000000",
        "00000000",
        -- code 0x49
        "00000000",
        "00000000",
        "00111100",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x4A
        "00000000",
        "00000000",
        "00001111",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x4B
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "01101100",
        "01101100",
        "01111000",
        "01111000",
        "01101100",
        "01101100",
        "01100110",
        "01100110",
        "01100110",
        "00000000",
        "00000000",
        -- code 0x4C
        "00000000",
        "00000000",
        "01111000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110010",
        "01111110",
        "00000000",
        "00000000",
        -- code 0x4D
        "00000000",
        "00000000",
        "01000010",
        "01100110",
        "01111110",
        "01111110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00000000",
        "00000000",
        -- code 0x4E
        "00000000",
        "00000000",
        "01100011",
        "01100011",
        "01110011",
        "01110011",
        "01101011",
        "01101011",
        "01100111",
        "01100111",
        "01100011",
        "01100011",
        "01100011",
        "01100011",
        "00000000",
        "00000000",
        -- code 0x4F
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x50
        "00000000",
        "00000000",
        "01111100",
        "00110110",
        "00110110",
        "00110110",
        "00110110",
        "00111100",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "01111000",
        "00000000",
        "00000000",
        -- code 0x51
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01101110",
        "01101110",
        "01101110",
        "00111100",
        "00001110",
        "00000000",
        -- code 0x52
        "00000000",
        "00000000",
        "01111110",
        "00110011",
        "00110011",
        "00110011",
        "00110011",
        "00111110",
        "00110110",
        "00110011",
        "00110011",
        "00110011",
        "00110011",
        "01111011",
        "00000000",
        "00000000",
        -- code 0x53
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "01100000",
        "00110000",
        "00011000",
        "00001100",
        "00000110",
        "00000110",
        "01100110",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x54
        "00000000",
        "00000000",
        "01111110",
        "01011010",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x55
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x56
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00111100",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        -- code 0x57
        "00000000",
        "00000000",
        "01100011",
        "01100011",
        "01100011",
        "01100011",
        "01100011",
        "01100011",
        "01100011",
        "01101011",
        "01101011",
        "01101011",
        "00111110",
        "00110110",
        "00000000",
        "00000000",
        -- code 0x58
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00111100",
        "00011000",
        "00011000",
        "00111100",
        "00111100",
        "01100110",
        "01100110",
        "01100110",
        "00000000",
        "00000000",
        -- code 0x59
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00111100",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x5A
        "00000000",
        "00000000",
        "01111110",
        "01000110",
        "00000110",
        "00001100",
        "00001100",
        "00011000",
        "00011000",
        "00110000",
        "00110000",
        "01100000",
        "01100010",
        "01111110",
        "00000000",
        "00000000",
        -- code 0x5B
        "00000000",
        "00111100",
        "00111100",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00111100",
        "00111100",
        "00000000",
        -- code 0x5C
        "00000000",
        "00000000",
        "01000000",
        "01100000",
        "01100000",
        "00110000",
        "00110000",
        "00011000",
        "00011000",
        "00001100",
        "00001100",
        "00000110",
        "00000110",
        "00000010",
        "00000000",
        "00000000",
        -- code 0x5D
        "00000000",
        "00111100",
        "00111100",
        "00001100",
        "00001100",
        "00001100",
        "00001100",
        "00001100",
        "00001100",
        "00001100",
        "00001100",
        "00001100",
        "00001100",
        "00111100",
        "00111100",
        "00000000",
        -- code 0x5E
        "00000000",
        "00000000",
        "00011000",
        "00111100",
        "01100110",
        "01000010",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x5F
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01111110",
        "00000000",
        -- code 0x60
        "00000000",
        "00100000",
        "00110000",
        "00110000",
        "00011000",
        "00011000",
        "00001000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x61
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "00000110",
        "00111110",
        "01100110",
        "01100110",
        "01101110",
        "00110111",
        "00000000",
        "00000000",
        -- code 0x62
        "00000000",
        "00000000",
        "01110000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00111100",
        "00110110",
        "00110110",
        "00110110",
        "00110110",
        "00110110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x63
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100000",
        "01100000",
        "01100000",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x64
        "00000000",
        "00000000",
        "00011100",
        "00001100",
        "00001100",
        "00001100",
        "00001100",
        "00111100",
        "01101100",
        "01101100",
        "01101100",
        "01101100",
        "01101100",
        "00110110",
        "00000000",
        "00000000",
        -- code 0x65
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "01111110",
        "01100000",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x66
        "00000000",
        "00000000",
        "00000000",
        "00011100",
        "00110110",
        "00110110",
        "00110000",
        "00110000",
        "01111000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "01111000",
        "00000000",
        "00000000",
        -- code 0x67
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111011",
        "01100110",
        "01100110",
        "01100110",
        "00111110",
        "00000110",
        "00000110",
        "01100110",
        "00111100",
        -- code 0x68
        "00000000",
        "00000000",
        "00000000",
        "01110000",
        "00110000",
        "00110000",
        "00110000",
        "00111100",
        "00110110",
        "00110110",
        "00110110",
        "00110110",
        "00110110",
        "01110110",
        "00000000",
        "00000000",
        -- code 0x69
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00000000",
        "00111000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x6A
        "00000000",
        "00000000",
        "00000000",
        "00000110",
        "00000110",
        "00000000",
        "00001110",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "00000110",
        "01100110",
        "01100110",
        "00111100",
        -- code 0x6B
        "00000000",
        "00000000",
        "01110000",
        "00110000",
        "00110000",
        "00110000",
        "00110011",
        "00110110",
        "00111100",
        "00111100",
        "00110110",
        "00110110",
        "00110011",
        "01110011",
        "00000000",
        "00000000",
        -- code 0x6C
        "00000000",
        "00000000",
        "00111000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x6D
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01110110",
        "01111111",
        "01101011",
        "01101011",
        "01101011",
        "01101011",
        "01101011",
        "00000000",
        "00000000",
        -- code 0x6E
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01101100",
        "00110110",
        "00110110",
        "00110110",
        "00110110",
        "00110110",
        "00110110",
        "00000000",
        "00000000",
        -- code 0x6F
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x70
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01011110",
        "00110011",
        "00110011",
        "00110011",
        "00110011",
        "00111110",
        "00110000",
        "00110000",
        "00110000",
        -- code 0x71
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111101",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111110",
        "00000110",
        "00000110",
        "00000110",
        -- code 0x72
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01011100",
        "00110110",
        "00110110",
        "00110000",
        "00110000",
        "00110000",
        "01111000",
        "00000000",
        "00000000",
        -- code 0x73
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "01100110",
        "00110000",
        "00011000",
        "00001100",
        "01100110",
        "00111100",
        "00000000",
        "00000000",
        -- code 0x74
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00010000",
        "00110000",
        "00110000",
        "01111000",
        "00110000",
        "00110000",
        "00110000",
        "00110000",
        "00110110",
        "00011100",
        "00000000",
        "00000000",
        -- code 0x75
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01101100",
        "01101100",
        "01101100",
        "01101100",
        "01101100",
        "01101100",
        "00111010",
        "00000000",
        "00000000",
        -- code 0x76
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111100",
        "00011000",
        "00000000",
        "00000000",
        -- code 0x77
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01100011",
        "01100011",
        "01100011",
        "01101011",
        "01101011",
        "00111110",
        "00110110",
        "00000000",
        "00000000",
        -- code 0x78
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01000010",
        "01100110",
        "00111100",
        "00011000",
        "00111100",
        "01100110",
        "01000010",
        "00000000",
        "00000000",
        -- code 0x79
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "01100110",
        "00111110",
        "00000110",
        "01000110",
        "00111100",
        -- code 0x7A
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01111110",
        "01000110",
        "00001100",
        "00011000",
        "00110000",
        "01100010",
        "01111110",
        "00000000",
        "00000000",
        -- code 0x7B
        "00000000",
        "01110000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00001110",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "01110000",
        "00000000",
        "00000000",
        -- code 0x7C
        "00000000",
        "00000000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00000000",
        "00000000",
        -- code 0x7D
        "00000000",
        "00001110",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "01110000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00011000",
        "00001110",
        "00000000",
        "00000000",
        -- code 0x7E
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00110000",
        "01011010",
        "00001100",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        -- code 0x7F
        "00000000",
        "01111110",
        "01000010",
        "01000010",
        "01000010",
        "01000010",
        "01000010",
        "01000010",
        "01000010",
        "01000010",
        "01000010",
        "01000010",
        "01000010",
        "01000010",
        "01111110",
        "00000000"
    );

begin

    process (clk) is
    begin

        if rising_edge(clk) then
            data <= ROM(to_integer(addr));
        end if;

    end process;

end architecture font_rom_arch;
